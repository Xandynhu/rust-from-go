module top_module(
    input logic clk,
    input logic rst_n,
    input logic [7:0] data_in,
    output logic [7:0] data_out,
    inout logic bidir_port,
    output logic [3:0] multi_bit_out,
    input logic [3:0] multi_bit_in
);

    // Instantiate module_with_ports
    module_with_ports module_inst(
        .clk(clk),
        .rst_n(rst_n),
        .data_in(data_in),
        .data_out(data_out),
        .bidir_port(bidir_port),
        .multi_bit_out(multi_bit_out),
        .multi_bit_in(multi_bit_in)
    );

endmodule
